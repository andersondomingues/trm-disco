module fetch(


);


endmodule